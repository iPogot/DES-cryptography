module key_generator #(parameter KEY_WIDTH = 48
)
(

);





    

endmodule